module Unified_Buffer #(
) (
);

endmodule

