module Accumulator_tb ();
endmodule
